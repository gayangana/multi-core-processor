module CID #( parameter cid)(
    output [15:0] data_out
);


assign  data_out = cid;
endmodule

